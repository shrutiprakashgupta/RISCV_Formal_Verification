module tb_top (

input        clk_i,
input        reset_i,
input [31:0] iaddr_o 
);

endmodule
